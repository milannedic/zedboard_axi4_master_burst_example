`timescale 1 ns / 1 ps

module axi_datamover_wrap
(

 input logic                 m_axi_mm2s_aclk,
 input logic                 m_axi_mm2s_aresetn,
 input logic                 m_axis_mm2s_cmdsts_aclk,
 input logic                 m_axis_mm2s_cmdsts_aresetn,
 input logic                 s_axis_mm2s_cmd_tvalid,
 output logic                s_axis_mm2s_cmd_tready,
 input logic [40+32-1: 0]    s_axis_mm2s_cmd_tdata,
 output logic                m_axis_mm2s_sts_tvalid,
 input logic                 m_axis_mm2s_sts_tready,
 output logic [7 : 0]        m_axis_mm2s_sts_tdata,
 output logic [0 : 0]        m_axis_mm2s_sts_tkeep,
 output logic                m_axis_mm2s_sts_tlast,
 output logic [4-1 : 0]      m_axi_mm2s_arid,
 output logic [32-1 : 0]     m_axi_mm2s_araddr,
 output logic [7 : 0]        m_axi_mm2s_arlen,
 output logic [2 : 0]        m_axi_mm2s_arsize,
 output logic [1 : 0]        m_axi_mm2s_arburst,
 output logic [2 : 0]        m_axi_mm2s_arprot,
 output logic [3 : 0]        m_axi_mm2s_arcache,
 output logic [3 : 0]        m_axi_mm2s_aruser,
 output logic                m_axi_mm2s_arvalid,
 input logic                 m_axi_mm2s_arready,
 input logic [64-1 : 0]      m_axi_mm2s_rdata,
 input logic [1 : 0]         m_axi_mm2s_rresp,
 input logic                 m_axi_mm2s_rlast,
 input logic                 m_axi_mm2s_rvalid,
 output logic                m_axi_mm2s_rready,
 output logic [64-1 : 0]     m_axis_mm2s_tdata,
 output logic [(64/8)-1 : 0] m_axis_mm2s_tkeep,
 output logic                m_axis_mm2s_tlast,
 output logic                m_axis_mm2s_tvalid,
 input logic                 m_axis_mm2s_tready,
 output logic                mm2s_err,
 input logic                 m_axi_s2mm_aclk,
 input logic                 m_axi_s2mm_aresetn,
 input logic                 m_axis_s2mm_cmdsts_awclk,
 input logic                 m_axis_s2mm_cmdsts_aresetn,
 input logic                 s_axis_s2mm_cmd_tvalid,
 output logic                s_axis_s2mm_cmd_tready,
 input logic [40+32-1 : 0]   s_axis_s2mm_cmd_tdata,
 output logic                m_axis_s2mm_sts_tvalid,
 input logic                 m_axis_s2mm_sts_tready,
 output logic [7 : 0]        m_axis_s2mm_sts_tdata,
 output logic [0 : 0]        m_axis_s2mm_sts_tkeep,
 output logic                m_axis_s2mm_sts_tlast,
 output logic [4-1 : 0]      m_axi_s2mm_awid,
 output logic [32-1 : 0]     m_axi_s2mm_awaddr,
 output logic [7 : 0]        m_axi_s2mm_awlen,
 output logic [2 : 0]        m_axi_s2mm_awsize,
 output logic [1 : 0]        m_axi_s2mm_awburst,
 output logic [2 : 0]        m_axi_s2mm_awprot,
 output logic [3 : 0]        m_axi_s2mm_awcache,
 output logic [3 : 0]        m_axi_s2mm_awuser,
 output logic                m_axi_s2mm_awvalid,
 input logic                 m_axi_s2mm_awready,
 output logic [64-1 : 0]     m_axi_s2mm_wdata,
 output logic [(64/8)-1 : 0] m_axi_s2mm_wstrb,
 output logic                m_axi_s2mm_wlast,
 output logic                m_axi_s2mm_wvalid,
 input logic                 m_axi_s2mm_wready,
 input logic [1 : 0]         m_axi_s2mm_bresp,
 input logic                 m_axi_s2mm_bvalid,
 output logic                m_axi_s2mm_bready,
 input logic [64-1 : 0]      s_axis_s2mm_tdata,
 input logic [(64/8)-1 : 0]  s_axis_s2mm_tkeep,
 input logic                 s_axis_s2mm_tlast,
 input logic                 s_axis_s2mm_tvalid,
 output logic                s_axis_s2mm_tready,
 output logic                s2mm_err
);

endmodule
